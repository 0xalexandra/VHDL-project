library verilog;
use verilog.vl_types.all;
entity problhma1_vlg_vec_tst is
end problhma1_vlg_vec_tst;
