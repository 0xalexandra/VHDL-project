library verilog;
use verilog.vl_types.all;
entity problhma3_vlg_vec_tst is
end problhma3_vlg_vec_tst;
