library verilog;
use verilog.vl_types.all;
entity problhma2_vlg_vec_tst is
end problhma2_vlg_vec_tst;
